
module clk_custom (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
